package q_8_34a_pkg;
    parameter data_size = 8;
    parameter r2_size = 4;
endpackage
