package q_8_34a_pkg;
    parameter data_size = 4;
    parameter r2_size = 2;
endpackage
