package state_pkg;
    typedef enum logic [1:0] {S_idle, S_1, S_2} state_t;
endpackage
