package q_8_37_pkg;
    parameter r2_size = 4;
    parameter data_size = 8;
    typedef enum logic {
        S_idle,
        S_running
    } state_t;
endpackage
