package q_8_29_rtl_pkg;
    typedef enum logic [2:0] {
        S_0, S_1, S_2, S_3, S_4, S_5, S_6, S_7
    } state_t;
endpackage
