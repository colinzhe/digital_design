package q_8_37c_pkg;
    parameter r2_size = 4;
    parameter data_size = 8;
endpackage
