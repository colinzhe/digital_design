package ex_8_8_pkg;
    parameter st_width = 3;
    typedef enum logic [st_width-1:0] {S0, S1, S2, S3} state_t;
    parameter r1_size = 8, r2_size = 4;
    //supply0 GND;
    //supply1 PWR;
endpackage
