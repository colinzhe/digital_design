module seven_seg (
    x,
    hexd
);
    input [3:0] x;
    output [6:0] hexd;
    
    assign hexd[0] = (~x[3] & x[2] & ~x[1] & ~x[0]) | (~x[3] & ~x[2] & ~x[1] & x[0])
        | (x[3] & x[2] & ~x[1] & x[0]) | (x[3] & ~x[2] & x[1] & x[0]);
        
    assign hexd[1] = (~x[3] & x[2] & ~x[1] & x[0]) | (x[2] & x[1] & ~x[0])
        | (x[3] & x[2] & ~x[0]) | (x[3] & x[2] & x[1]) | (x[3] & x[1] & x[0]);
        
    assign hexd[2] = (~x[3] & ~x[2] & x[1] & ~x[0]) | (x[3] & x[2] & ~x[1] & ~x[0])
        | (x[3] & x[2] & x[1]);
        
    assign hexd[3] = (~x[3] & ~x[2] & ~x[1] & x[0]) | (~x[3] & x[2] & ~x[1] & ~x[0])
        | (x[2] & x[1] & x[0]) | (x[3] & ~x[2] & x[1] & ~x[0]);
        
    assign hexd[4] = (~x[2] & ~x[1] & x[0]) | (~x[3] & x[0]) | (~x[3] & x[2] & ~x[1]);
    
    assign hexd[5] = (~x[3] & ~x[2] & x[0]) | (~x[3] & ~x[2] & x[1]) | (~x[3] & x[1] & x[0])
        | (x[3] & x[2] & ~x[1] & x[0]);
        
    assign hexd[6] = (~x[3] & ~x[2] & ~x[1]) | (~x[3] & x[2] & x[1] & x[0])
        | (x[3] & x[2] & ~x[1] & ~x[0]);
endmodule
