package q_8_7_pkg;
    parameter st_width = 2;
    typedef enum logic [st_width-1:0] {S_idle, S_1, S_2} state_t;
endpackage;
