package q_8_8_pkg;
    parameter st_width = 2;
    typedef enum logic [st_width-1:0] {
        S_idle, S_1
    } state_t;
endpackage
