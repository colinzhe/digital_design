package ex_8_8_pkg;
    enum logic [1:0] {S0, S1, S2, S3};
    parameter r1_size = 8, r2_size = 4;
    supply0 GND;
    supply1 PWR;
endpackage
