package q_8_28_pkg;
    parameter dp_width = 5;
    parameter bc_size = 3;
    parameter st_width = 3;
endpackage
