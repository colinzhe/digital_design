package q_8_34b_pkg;
    typedef enum logic [1:0] {
        S_idle,
        S_1,
        S_2,
        S_3
    } state_t;
endpackage
