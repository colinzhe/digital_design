package q_8_42_pkg;
    parameter data_size = 8;
    parameter r2_size = 4;
    typedef enum logic {
        S_idle,
        S_count
    } state_t;
endpackage
