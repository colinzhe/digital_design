package q_8_41_pkg;
    typedef enum logic [1:0] {
        S_idle,
        S_1,
        S_full,
        S_wait
    } state_t;
endpackage
