package mul_u64_pkg;
    typedef enum logic [2:0] {
        s_mp_0,
        s_mp_1,
        s_mp_2,
        s_mp_3,
        s_mp_final
    } mult_pass_t;