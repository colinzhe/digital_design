package q_8_39_pkg;
    parameter data_width = 4;
endpackage
